`define PKT_PREAMBLE    8'hCA
`define PKT_COMMAND_CPU_WRITE 4'h1
`define PKT_COMMAND_CPU_READ  4'h2
`define PKT_COMMAND_DAQ_WRITE 4'h3
`define PKT_COMMAND_DAQ_READ  4'h4
