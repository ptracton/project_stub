//                              -*- Mode: Verilog -*-
// Filename        : wb_dsp_includes.vh
// Description     : Include file for WB DSP Testing
// Author          : Philip Tracton
// Created On      : Wed Dec  2 13:38:15 2015
// Last Modified By: Philip Tracton
// Last Modified On: Wed Dec  2 13:38:15 2015
// Update Count    : 0
// Status          : Unknown, Use with caution!



`define WB_RAM0 19'h4_0000
`define WB_RAM1 19'h4_2000
`define WB_RAM2 19'h4_4000
`define WB_RAM3 19'h4_6000


`define WB_FULL_WORD       4'hF
`define WB_UPPER_HALF_WORD 4'hC
`define WB_LOWER_HALF_WORD 4'h3
`define WB_BYTE_0          4'h1
`define WB_BYTE_1          4'h2
`define WB_BYTE_2          4'h4
`define WB_BYTE_3          4'h8
